//for dot matrix
//Frequency Divider: Transfer the frequency to 10000 Hz (instead of 50MHz)
`define TimeExpire 32'd2500

module FrequencyDivider2(clk, rst, div_clk);
input clk, rst;
output div_clk;

reg div_clk;
reg [31:0] count;

always @(posedge clk)
begin
	if(!rst) //low Sycn reset
	begin
		count <= 32'd0;
		div_clk <= 32'd0;
	end
	
	else
	begin
		if(count == `TimeExpire)
		begin
			count <= 32'd0;
			div_clk <= ~div_clk;
			
		end
		
		else
		begin
			count <= count + 32'd1;	
		end 
		
	end


end

endmodule